
module unsaved (
	clk_clk,
	reset_reset_n,
	pll_0_sdram_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		pll_0_sdram_clk;
endmodule
