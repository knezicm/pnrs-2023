-- soc_system.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                           : in    std_logic                     := '0';             --                     clk.clk
		hps_0_ddr_mem_a                   : out   std_logic_vector(14 downto 0);                    --               hps_0_ddr.mem_a
		hps_0_ddr_mem_ba                  : out   std_logic_vector(2 downto 0);                     --                        .mem_ba
		hps_0_ddr_mem_ck                  : out   std_logic;                                        --                        .mem_ck
		hps_0_ddr_mem_ck_n                : out   std_logic;                                        --                        .mem_ck_n
		hps_0_ddr_mem_cke                 : out   std_logic;                                        --                        .mem_cke
		hps_0_ddr_mem_cs_n                : out   std_logic;                                        --                        .mem_cs_n
		hps_0_ddr_mem_ras_n               : out   std_logic;                                        --                        .mem_ras_n
		hps_0_ddr_mem_cas_n               : out   std_logic;                                        --                        .mem_cas_n
		hps_0_ddr_mem_we_n                : out   std_logic;                                        --                        .mem_we_n
		hps_0_ddr_mem_reset_n             : out   std_logic;                                        --                        .mem_reset_n
		hps_0_ddr_mem_dq                  : inout std_logic_vector(31 downto 0) := (others => '0'); --                        .mem_dq
		hps_0_ddr_mem_dqs                 : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs
		hps_0_ddr_mem_dqs_n               : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs_n
		hps_0_ddr_mem_odt                 : out   std_logic;                                        --                        .mem_odt
		hps_0_ddr_mem_dm                  : out   std_logic_vector(3 downto 0);                     --                        .mem_dm
		hps_0_ddr_oct_rzqin               : in    std_logic                     := '0';             --                        .oct_rzqin
		hps_0_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --                hps_0_io.hps_io_emac1_inst_TX_CLK
		hps_0_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD0
		hps_0_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD1
		hps_0_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD2
		hps_0_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD3
		hps_0_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD0
		hps_0_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                        .hps_io_emac1_inst_MDIO
		hps_0_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                        .hps_io_emac1_inst_MDC
		hps_0_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CTL
		hps_0_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                        .hps_io_emac1_inst_TX_CTL
		hps_0_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CLK
		hps_0_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD1
		hps_0_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD2
		hps_0_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD3
		hps_0_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_CMD
		hps_0_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D0
		hps_0_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D1
		hps_0_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                        .hps_io_sdio_inst_CLK
		hps_0_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D2
		hps_0_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D3
		hps_0_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                        .hps_io_uart0_inst_RX
		hps_0_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                        .hps_io_uart0_inst_TX
		hps_0_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO35
		hps_0_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO53
		hps_0_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO54
		pll_0_sdram_clk                   : out   std_logic;                                        --             pll_0_sdram.clk
		reset_reset_n                     : in    std_logic                     := '0';             --                   reset.reset_n
		sdram_controller_0_wire_addr      : out   std_logic_vector(12 downto 0);                    -- sdram_controller_0_wire.addr
		sdram_controller_0_wire_ba        : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_controller_0_wire_cas_n     : out   std_logic;                                        --                        .cas_n
		sdram_controller_0_wire_cke       : out   std_logic;                                        --                        .cke
		sdram_controller_0_wire_cs_n      : out   std_logic;                                        --                        .cs_n
		sdram_controller_0_wire_dq        : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_controller_0_wire_dqm       : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_controller_0_wire_ras_n     : out   std_logic;                                        --                        .ras_n
		sdram_controller_0_wire_we_n      : out   std_logic                                         --                        .we_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_finished_mutex is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component soc_system_finished_mutex;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component soc_system_hps_0;

	component soc_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart_0;

	component soc_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_pll_0;

	component soc_system_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component soc_system_sdram_controller_0;

	component soc_system_smoker_with_matches is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_smoker_with_matches;

	component soc_system_smoker_with_paper is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_smoker_with_paper;

	component soc_system_smoker_with_tobacco is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_smoker_with_tobacco;

	component soc_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid;

	component soc_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_timer_0;

	component soc_system_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			pll_0_outclk0_clk                                                   : in  std_logic                     := 'X';             -- clk
			pll_0_outclk1_clk                                                   : in  std_logic                     := 'X';             -- clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			sdram_controller_0_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			smoker_with_matches_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			smoker_with_paper_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			smoker_with_tobacco_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			timer_1_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			timer_2_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			tobacco_mutex_reset_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			smoker_with_matches_data_master_address                             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_matches_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			smoker_with_matches_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			smoker_with_matches_data_master_read                                : in  std_logic                     := 'X';             -- read
			smoker_with_matches_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			smoker_with_matches_data_master_write                               : in  std_logic                     := 'X';             -- write
			smoker_with_matches_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			smoker_with_matches_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			smoker_with_matches_instruction_master_address                      : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_matches_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			smoker_with_matches_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			smoker_with_matches_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			smoker_with_paper_data_master_address                               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_paper_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			smoker_with_paper_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			smoker_with_paper_data_master_read                                  : in  std_logic                     := 'X';             -- read
			smoker_with_paper_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			smoker_with_paper_data_master_write                                 : in  std_logic                     := 'X';             -- write
			smoker_with_paper_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			smoker_with_paper_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			smoker_with_paper_instruction_master_address                        : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_paper_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			smoker_with_paper_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			smoker_with_paper_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			smoker_with_tobacco_data_master_address                             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_tobacco_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			smoker_with_tobacco_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			smoker_with_tobacco_data_master_read                                : in  std_logic                     := 'X';             -- read
			smoker_with_tobacco_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			smoker_with_tobacco_data_master_write                               : in  std_logic                     := 'X';             -- write
			smoker_with_tobacco_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			smoker_with_tobacco_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			smoker_with_tobacco_instruction_master_address                      : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			smoker_with_tobacco_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			smoker_with_tobacco_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			smoker_with_tobacco_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			finished_mutex_s1_address                                           : out std_logic_vector(0 downto 0);                     -- address
			finished_mutex_s1_write                                             : out std_logic;                                        -- write
			finished_mutex_s1_read                                              : out std_logic;                                        -- read
			finished_mutex_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			finished_mutex_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			finished_mutex_s1_chipselect                                        : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                                 : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                                  : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                            : out std_logic;                                        -- chipselect
			matches_mutex_s1_address                                            : out std_logic_vector(0 downto 0);                     -- address
			matches_mutex_s1_write                                              : out std_logic;                                        -- write
			matches_mutex_s1_read                                               : out std_logic;                                        -- read
			matches_mutex_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			matches_mutex_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			matches_mutex_s1_chipselect                                         : out std_logic;                                        -- chipselect
			paper_mutex_s1_address                                              : out std_logic_vector(0 downto 0);                     -- address
			paper_mutex_s1_write                                                : out std_logic;                                        -- write
			paper_mutex_s1_read                                                 : out std_logic;                                        -- read
			paper_mutex_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			paper_mutex_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			paper_mutex_s1_chipselect                                           : out std_logic;                                        -- chipselect
			sdram_controller_0_s1_address                                       : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_0_s1_write                                         : out std_logic;                                        -- write
			sdram_controller_0_s1_read                                          : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable                                    : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid                                 : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest                                   : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect                                    : out std_logic;                                        -- chipselect
			smoker_with_matches_debug_mem_slave_address                         : out std_logic_vector(8 downto 0);                     -- address
			smoker_with_matches_debug_mem_slave_write                           : out std_logic;                                        -- write
			smoker_with_matches_debug_mem_slave_read                            : out std_logic;                                        -- read
			smoker_with_matches_debug_mem_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			smoker_with_matches_debug_mem_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			smoker_with_matches_debug_mem_slave_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			smoker_with_matches_debug_mem_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			smoker_with_matches_debug_mem_slave_debugaccess                     : out std_logic;                                        -- debugaccess
			smoker_with_paper_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			smoker_with_paper_debug_mem_slave_write                             : out std_logic;                                        -- write
			smoker_with_paper_debug_mem_slave_read                              : out std_logic;                                        -- read
			smoker_with_paper_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			smoker_with_paper_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			smoker_with_paper_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			smoker_with_paper_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			smoker_with_paper_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			smoker_with_tobacco_debug_mem_slave_address                         : out std_logic_vector(8 downto 0);                     -- address
			smoker_with_tobacco_debug_mem_slave_write                           : out std_logic;                                        -- write
			smoker_with_tobacco_debug_mem_slave_read                            : out std_logic;                                        -- read
			smoker_with_tobacco_debug_mem_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			smoker_with_tobacco_debug_mem_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			smoker_with_tobacco_debug_mem_slave_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			smoker_with_tobacco_debug_mem_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			smoker_with_tobacco_debug_mem_slave_debugaccess                     : out std_logic;                                        -- debugaccess
			sysid_control_slave_address                                         : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                                    : out std_logic;                                        -- write
			timer_0_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                               : out std_logic;                                        -- chipselect
			timer_1_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                                    : out std_logic;                                        -- write
			timer_1_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                                               : out std_logic;                                        -- chipselect
			timer_2_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			timer_2_s1_write                                                    : out std_logic;                                        -- write
			timer_2_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_2_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_2_s1_chipselect                                               : out std_logic;                                        -- chipselect
			tobacco_mutex_s1_address                                            : out std_logic_vector(0 downto 0);                     -- address
			tobacco_mutex_s1_write                                              : out std_logic;                                        -- write
			tobacco_mutex_s1_read                                               : out std_logic;                                        -- read
			tobacco_mutex_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tobacco_mutex_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			tobacco_mutex_s1_chipselect                                         : out std_logic                                         -- chipselect
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			reset_in3      : in  std_logic := 'X'; -- reset_in3.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	component soc_system_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_003;

	component soc_system_rst_controller_005 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_005;

	component soc_system_rst_controller_006 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_006;

	signal pll_0_outclk0_clk                                                 : std_logic;                     -- pll_0:outclk_0 -> [finished_mutex:clk, hps_0:h2f_lw_axi_clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, jtag_uart_0:clk, matches_mutex:clk, mm_interconnect_0:pll_0_outclk0_clk, paper_mutex:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_004:clk, rst_controller_005:clk, rst_controller_006:clk, rst_controller_007:clk, rst_controller_008:clk, smoker_with_paper:clk, smoker_with_tobacco:clk, sysid:clock, timer_0:clk, timer_1:clk, timer_2:clk, tobacco_mutex:clk]
	signal pll_0_outclk1_clk                                                 : std_logic;                     -- pll_0:outclk_1 -> [mm_interconnect_0:pll_0_outclk1_clk, rst_controller_002:clk, sdram_controller_0:clk]
	signal smoker_with_tobacco_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_tobacco_data_master_readdata -> smoker_with_tobacco:d_readdata
	signal smoker_with_tobacco_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:smoker_with_tobacco_data_master_waitrequest -> smoker_with_tobacco:d_waitrequest
	signal smoker_with_tobacco_data_master_debugaccess                       : std_logic;                     -- smoker_with_tobacco:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:smoker_with_tobacco_data_master_debugaccess
	signal smoker_with_tobacco_data_master_address                           : std_logic_vector(26 downto 0); -- smoker_with_tobacco:d_address -> mm_interconnect_0:smoker_with_tobacco_data_master_address
	signal smoker_with_tobacco_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- smoker_with_tobacco:d_byteenable -> mm_interconnect_0:smoker_with_tobacco_data_master_byteenable
	signal smoker_with_tobacco_data_master_read                              : std_logic;                     -- smoker_with_tobacco:d_read -> mm_interconnect_0:smoker_with_tobacco_data_master_read
	signal smoker_with_tobacco_data_master_write                             : std_logic;                     -- smoker_with_tobacco:d_write -> mm_interconnect_0:smoker_with_tobacco_data_master_write
	signal smoker_with_tobacco_data_master_writedata                         : std_logic_vector(31 downto 0); -- smoker_with_tobacco:d_writedata -> mm_interconnect_0:smoker_with_tobacco_data_master_writedata
	signal smoker_with_paper_data_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_paper_data_master_readdata -> smoker_with_paper:d_readdata
	signal smoker_with_paper_data_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:smoker_with_paper_data_master_waitrequest -> smoker_with_paper:d_waitrequest
	signal smoker_with_paper_data_master_debugaccess                         : std_logic;                     -- smoker_with_paper:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:smoker_with_paper_data_master_debugaccess
	signal smoker_with_paper_data_master_address                             : std_logic_vector(26 downto 0); -- smoker_with_paper:d_address -> mm_interconnect_0:smoker_with_paper_data_master_address
	signal smoker_with_paper_data_master_byteenable                          : std_logic_vector(3 downto 0);  -- smoker_with_paper:d_byteenable -> mm_interconnect_0:smoker_with_paper_data_master_byteenable
	signal smoker_with_paper_data_master_read                                : std_logic;                     -- smoker_with_paper:d_read -> mm_interconnect_0:smoker_with_paper_data_master_read
	signal smoker_with_paper_data_master_write                               : std_logic;                     -- smoker_with_paper:d_write -> mm_interconnect_0:smoker_with_paper_data_master_write
	signal smoker_with_paper_data_master_writedata                           : std_logic_vector(31 downto 0); -- smoker_with_paper:d_writedata -> mm_interconnect_0:smoker_with_paper_data_master_writedata
	signal smoker_with_matches_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_matches_data_master_readdata -> smoker_with_matches:d_readdata
	signal smoker_with_matches_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:smoker_with_matches_data_master_waitrequest -> smoker_with_matches:d_waitrequest
	signal smoker_with_matches_data_master_debugaccess                       : std_logic;                     -- smoker_with_matches:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:smoker_with_matches_data_master_debugaccess
	signal smoker_with_matches_data_master_address                           : std_logic_vector(26 downto 0); -- smoker_with_matches:d_address -> mm_interconnect_0:smoker_with_matches_data_master_address
	signal smoker_with_matches_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- smoker_with_matches:d_byteenable -> mm_interconnect_0:smoker_with_matches_data_master_byteenable
	signal smoker_with_matches_data_master_read                              : std_logic;                     -- smoker_with_matches:d_read -> mm_interconnect_0:smoker_with_matches_data_master_read
	signal smoker_with_matches_data_master_write                             : std_logic;                     -- smoker_with_matches:d_write -> mm_interconnect_0:smoker_with_matches_data_master_write
	signal smoker_with_matches_data_master_writedata                         : std_logic_vector(31 downto 0); -- smoker_with_matches:d_writedata -> mm_interconnect_0:smoker_with_matches_data_master_writedata
	signal smoker_with_tobacco_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_tobacco_instruction_master_readdata -> smoker_with_tobacco:i_readdata
	signal smoker_with_tobacco_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:smoker_with_tobacco_instruction_master_waitrequest -> smoker_with_tobacco:i_waitrequest
	signal smoker_with_tobacco_instruction_master_address                    : std_logic_vector(26 downto 0); -- smoker_with_tobacco:i_address -> mm_interconnect_0:smoker_with_tobacco_instruction_master_address
	signal smoker_with_tobacco_instruction_master_read                       : std_logic;                     -- smoker_with_tobacco:i_read -> mm_interconnect_0:smoker_with_tobacco_instruction_master_read
	signal smoker_with_paper_instruction_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_paper_instruction_master_readdata -> smoker_with_paper:i_readdata
	signal smoker_with_paper_instruction_master_waitrequest                  : std_logic;                     -- mm_interconnect_0:smoker_with_paper_instruction_master_waitrequest -> smoker_with_paper:i_waitrequest
	signal smoker_with_paper_instruction_master_address                      : std_logic_vector(26 downto 0); -- smoker_with_paper:i_address -> mm_interconnect_0:smoker_with_paper_instruction_master_address
	signal smoker_with_paper_instruction_master_read                         : std_logic;                     -- smoker_with_paper:i_read -> mm_interconnect_0:smoker_with_paper_instruction_master_read
	signal smoker_with_matches_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_matches_instruction_master_readdata -> smoker_with_matches:i_readdata
	signal smoker_with_matches_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:smoker_with_matches_instruction_master_waitrequest -> smoker_with_matches:i_waitrequest
	signal smoker_with_matches_instruction_master_address                    : std_logic_vector(26 downto 0); -- smoker_with_matches:i_address -> mm_interconnect_0:smoker_with_matches_instruction_master_address
	signal smoker_with_matches_instruction_master_read                       : std_logic;                     -- smoker_with_matches:i_read -> mm_interconnect_0:smoker_with_matches_instruction_master_read
	signal hps_0_h2f_lw_axi_master_awburst                                   : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                    : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                       : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                    : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                       : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                                   : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                    : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                    : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                     : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                                   : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                                   : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                      : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                    : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                    : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                    : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                                   : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                                   : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                                   : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                    : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                     : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                     : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                      : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                       : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                    : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                                   : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                    : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect        : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata          : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest       : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read              : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write             : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                    : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- smoker_with_tobacco:debug_mem_slave_readdata -> mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_readdata
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_waitrequest : std_logic;                     -- smoker_with_tobacco:debug_mem_slave_waitrequest -> mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_waitrequest
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_debugaccess -> smoker_with_tobacco:debug_mem_slave_debugaccess
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_address -> smoker_with_tobacco:debug_mem_slave_address
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_read -> smoker_with_tobacco:debug_mem_slave_read
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_byteenable -> smoker_with_tobacco:debug_mem_slave_byteenable
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_write -> smoker_with_tobacco:debug_mem_slave_write
	signal mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_tobacco_debug_mem_slave_writedata -> smoker_with_tobacco:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_tobacco_mutex_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:tobacco_mutex_s1_chipselect -> tobacco_mutex:chipselect
	signal mm_interconnect_0_tobacco_mutex_s1_readdata                       : std_logic_vector(31 downto 0); -- tobacco_mutex:data_to_cpu -> mm_interconnect_0:tobacco_mutex_s1_readdata
	signal mm_interconnect_0_tobacco_mutex_s1_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:tobacco_mutex_s1_address -> tobacco_mutex:address
	signal mm_interconnect_0_tobacco_mutex_s1_read                           : std_logic;                     -- mm_interconnect_0:tobacco_mutex_s1_read -> tobacco_mutex:read
	signal mm_interconnect_0_tobacco_mutex_s1_write                          : std_logic;                     -- mm_interconnect_0:tobacco_mutex_s1_write -> tobacco_mutex:write
	signal mm_interconnect_0_tobacco_mutex_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:tobacco_mutex_s1_writedata -> tobacco_mutex:data_from_cpu
	signal mm_interconnect_0_paper_mutex_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:paper_mutex_s1_chipselect -> paper_mutex:chipselect
	signal mm_interconnect_0_paper_mutex_s1_readdata                         : std_logic_vector(31 downto 0); -- paper_mutex:data_to_cpu -> mm_interconnect_0:paper_mutex_s1_readdata
	signal mm_interconnect_0_paper_mutex_s1_address                          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:paper_mutex_s1_address -> paper_mutex:address
	signal mm_interconnect_0_paper_mutex_s1_read                             : std_logic;                     -- mm_interconnect_0:paper_mutex_s1_read -> paper_mutex:read
	signal mm_interconnect_0_paper_mutex_s1_write                            : std_logic;                     -- mm_interconnect_0:paper_mutex_s1_write -> paper_mutex:write
	signal mm_interconnect_0_paper_mutex_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:paper_mutex_s1_writedata -> paper_mutex:data_from_cpu
	signal mm_interconnect_0_matches_mutex_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:matches_mutex_s1_chipselect -> matches_mutex:chipselect
	signal mm_interconnect_0_matches_mutex_s1_readdata                       : std_logic_vector(31 downto 0); -- matches_mutex:data_to_cpu -> mm_interconnect_0:matches_mutex_s1_readdata
	signal mm_interconnect_0_matches_mutex_s1_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:matches_mutex_s1_address -> matches_mutex:address
	signal mm_interconnect_0_matches_mutex_s1_read                           : std_logic;                     -- mm_interconnect_0:matches_mutex_s1_read -> matches_mutex:read
	signal mm_interconnect_0_matches_mutex_s1_write                          : std_logic;                     -- mm_interconnect_0:matches_mutex_s1_write -> matches_mutex:write
	signal mm_interconnect_0_matches_mutex_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:matches_mutex_s1_writedata -> matches_mutex:data_from_cpu
	signal mm_interconnect_0_finished_mutex_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:finished_mutex_s1_chipselect -> finished_mutex:chipselect
	signal mm_interconnect_0_finished_mutex_s1_readdata                      : std_logic_vector(31 downto 0); -- finished_mutex:data_to_cpu -> mm_interconnect_0:finished_mutex_s1_readdata
	signal mm_interconnect_0_finished_mutex_s1_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:finished_mutex_s1_address -> finished_mutex:address
	signal mm_interconnect_0_finished_mutex_s1_read                          : std_logic;                     -- mm_interconnect_0:finished_mutex_s1_read -> finished_mutex:read
	signal mm_interconnect_0_finished_mutex_s1_write                         : std_logic;                     -- mm_interconnect_0:finished_mutex_s1_write -> finished_mutex:write
	signal mm_interconnect_0_finished_mutex_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:finished_mutex_s1_writedata -> finished_mutex:data_from_cpu
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata                  : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest               : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address                   : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                      : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid             : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                     : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- smoker_with_matches:debug_mem_slave_readdata -> mm_interconnect_0:smoker_with_matches_debug_mem_slave_readdata
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_waitrequest : std_logic;                     -- smoker_with_matches:debug_mem_slave_waitrequest -> mm_interconnect_0:smoker_with_matches_debug_mem_slave_waitrequest
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_debugaccess -> smoker_with_matches:debug_mem_slave_debugaccess
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_address -> smoker_with_matches:debug_mem_slave_address
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_read -> smoker_with_matches:debug_mem_slave_read
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_byteenable -> smoker_with_matches:debug_mem_slave_byteenable
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_write -> smoker_with_matches:debug_mem_slave_write
	signal mm_interconnect_0_smoker_with_matches_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_matches_debug_mem_slave_writedata -> smoker_with_matches:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_2_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	signal mm_interconnect_0_timer_2_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	signal mm_interconnect_0_timer_2_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_2_s1_address -> timer_2:address
	signal mm_interconnect_0_timer_2_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_2_s1_write -> mm_interconnect_0_timer_2_s1_write:in
	signal mm_interconnect_0_timer_2_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_readdata      : std_logic_vector(31 downto 0); -- smoker_with_paper:debug_mem_slave_readdata -> mm_interconnect_0:smoker_with_paper_debug_mem_slave_readdata
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_waitrequest   : std_logic;                     -- smoker_with_paper:debug_mem_slave_waitrequest -> mm_interconnect_0:smoker_with_paper_debug_mem_slave_waitrequest
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_debugaccess   : std_logic;                     -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_debugaccess -> smoker_with_paper:debug_mem_slave_debugaccess
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_address       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_address -> smoker_with_paper:debug_mem_slave_address
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_read          : std_logic;                     -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_read -> smoker_with_paper:debug_mem_slave_read
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_byteenable -> smoker_with_paper:debug_mem_slave_byteenable
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_write         : std_logic;                     -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_write -> smoker_with_paper:debug_mem_slave_write
	signal mm_interconnect_0_smoker_with_paper_debug_mem_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:smoker_with_paper_debug_mem_slave_writedata -> smoker_with_paper:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal smoker_with_matches_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> smoker_with_matches:irq
	signal irq_mapper_001_receiver0_irq                                      : std_logic;                     -- timer_1:irq -> irq_mapper_001:receiver0_irq
	signal smoker_with_paper_irq_irq                                         : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> smoker_with_paper:irq
	signal irq_mapper_002_receiver1_irq                                      : std_logic;                     -- timer_0:irq -> irq_mapper_002:receiver1_irq
	signal smoker_with_tobacco_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> smoker_with_tobacco:irq
	signal irq_mapper_receiver0_irq                                          : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                     : std_logic_vector(0 downto 0);  -- timer_2:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                          : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_001_receiver1_irq                                      : std_logic;                     -- jtag_uart_0:av_irq -> [irq_mapper_001:receiver1_irq, irq_mapper_002:receiver0_irq, irq_synchronizer_001:receiver_irq]
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:tobacco_mutex_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal smoker_with_tobacco_debug_reset_request_reset                     : std_logic;                     -- smoker_with_tobacco:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_005:reset_in1]
	signal smoker_with_paper_debug_reset_request_reset                       : std_logic;                     -- smoker_with_paper:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_006:reset_in1]
	signal rst_controller_001_reset_out_reset                                : std_logic;                     -- rst_controller_001:reset_out -> [irq_synchronizer_001:receiver_reset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal smoker_with_matches_debug_reset_request_reset                     : std_logic;                     -- smoker_with_matches:debug_reset_request -> [rst_controller_001:reset_in3, rst_controller_007:reset_in1]
	signal rst_controller_002_reset_out_reset                                : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:sdram_controller_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                                : std_logic;                     -- rst_controller_003:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:smoker_with_matches_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_003_reset_out_reset_req                            : std_logic;                     -- rst_controller_003:reset_req -> [rst_translator:reset_req_in, smoker_with_matches:reset_req]
	signal rst_controller_004_reset_out_reset                                : std_logic;                     -- rst_controller_004:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:smoker_with_paper_reset_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in]
	signal rst_controller_004_reset_out_reset_req                            : std_logic;                     -- rst_controller_004:reset_req -> [rst_translator_001:reset_req_in, smoker_with_paper:reset_req]
	signal rst_controller_005_reset_out_reset                                : std_logic;                     -- rst_controller_005:reset_out -> [irq_mapper_002:reset, mm_interconnect_0:smoker_with_tobacco_reset_reset_bridge_in_reset_reset, rst_controller_005_reset_out_reset:in, rst_translator_002:in_reset]
	signal rst_controller_005_reset_out_reset_req                            : std_logic;                     -- rst_controller_005:reset_req -> [rst_translator_002:reset_req_in, smoker_with_tobacco:reset_req]
	signal rst_controller_006_reset_out_reset                                : std_logic;                     -- rst_controller_006:reset_out -> [mm_interconnect_0:timer_1_reset_reset_bridge_in_reset_reset, rst_controller_006_reset_out_reset:in]
	signal rst_controller_007_reset_out_reset                                : std_logic;                     -- rst_controller_007:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:timer_2_reset_reset_bridge_in_reset_reset, rst_controller_007_reset_out_reset:in]
	signal rst_controller_008_reset_out_reset                                : std_logic;                     -- rst_controller_008:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal hps_0_h2f_reset_reset                                             : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                           : std_logic;                     -- reset_reset_n:inv -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0, rst_controller_007:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv            : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv      : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal mm_interconnect_0_timer_2_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_2_s1_write:inv -> timer_2:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [finished_mutex:reset_n, matches_mutex:reset_n, paper_mutex:reset_n, tobacco_mutex:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart_0:rst_n, sysid:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> sdram_controller_0:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> smoker_with_matches:reset_n
	signal rst_controller_004_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> smoker_with_paper:reset_n
	signal rst_controller_005_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_005_reset_out_reset:inv -> [smoker_with_tobacco:reset_n, timer_0:reset_n]
	signal rst_controller_006_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_006_reset_out_reset:inv -> timer_1:reset_n
	signal rst_controller_007_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_007_reset_out_reset:inv -> timer_2:reset_n
	signal hps_0_h2f_reset_reset_ports_inv                                   : std_logic;                     -- hps_0_h2f_reset_reset:inv -> rst_controller_008:reset_in0

begin

	finished_mutex : component soc_system_finished_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,       -- reset.reset_n
			clk           => pll_0_outclk0_clk,                              --   clk.clk
			chipselect    => mm_interconnect_0_finished_mutex_s1_chipselect, --    s1.chipselect
			data_from_cpu => mm_interconnect_0_finished_mutex_s1_writedata,  --      .writedata
			read          => mm_interconnect_0_finished_mutex_s1_read,       --      .read
			write         => mm_interconnect_0_finished_mutex_s1_write,      --      .write
			data_to_cpu   => mm_interconnect_0_finished_mutex_s1_readdata,   --      .readdata
			address       => mm_interconnect_0_finished_mutex_s1_address(0)  --      .address
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => hps_0_ddr_mem_a,                   --            memory.mem_a
			mem_ba                   => hps_0_ddr_mem_ba,                  --                  .mem_ba
			mem_ck                   => hps_0_ddr_mem_ck,                  --                  .mem_ck
			mem_ck_n                 => hps_0_ddr_mem_ck_n,                --                  .mem_ck_n
			mem_cke                  => hps_0_ddr_mem_cke,                 --                  .mem_cke
			mem_cs_n                 => hps_0_ddr_mem_cs_n,                --                  .mem_cs_n
			mem_ras_n                => hps_0_ddr_mem_ras_n,               --                  .mem_ras_n
			mem_cas_n                => hps_0_ddr_mem_cas_n,               --                  .mem_cas_n
			mem_we_n                 => hps_0_ddr_mem_we_n,                --                  .mem_we_n
			mem_reset_n              => hps_0_ddr_mem_reset_n,             --                  .mem_reset_n
			mem_dq                   => hps_0_ddr_mem_dq,                  --                  .mem_dq
			mem_dqs                  => hps_0_ddr_mem_dqs,                 --                  .mem_dqs
			mem_dqs_n                => hps_0_ddr_mem_dqs_n,               --                  .mem_dqs_n
			mem_odt                  => hps_0_ddr_mem_odt,                 --                  .mem_odt
			mem_dm                   => hps_0_ddr_mem_dm,                  --                  .mem_dm
			oct_rzqin                => hps_0_ddr_oct_rzqin,               --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_io_hps_io_emac1_inst_TX_CLK, --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_io_hps_io_emac1_inst_TXD0,   --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_io_hps_io_emac1_inst_TXD1,   --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_io_hps_io_emac1_inst_TXD2,   --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_io_hps_io_emac1_inst_TXD3,   --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_io_hps_io_emac1_inst_RXD0,   --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_io_hps_io_emac1_inst_MDIO,   --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_io_hps_io_emac1_inst_MDC,    --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_io_hps_io_emac1_inst_RX_CTL, --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_io_hps_io_emac1_inst_TX_CTL, --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_io_hps_io_emac1_inst_RX_CLK, --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_io_hps_io_emac1_inst_RXD1,   --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_io_hps_io_emac1_inst_RXD2,   --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_io_hps_io_emac1_inst_RXD3,   --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_io_hps_io_sdio_inst_CMD,     --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_io_hps_io_sdio_inst_D0,      --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_io_hps_io_sdio_inst_D1,      --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_io_hps_io_sdio_inst_CLK,     --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_io_hps_io_sdio_inst_D2,      --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_io_hps_io_sdio_inst_D3,      --                  .hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     => hps_0_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO35  => hps_0_io_hps_io_gpio_inst_GPIO35,  --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO53  => hps_0_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_io_hps_io_gpio_inst_GPIO54,  --                  .hps_io_gpio_inst_GPIO54
			h2f_rst_n                => hps_0_h2f_reset_reset,             --         h2f_reset.reset_n
			h2f_lw_axi_clk           => pll_0_outclk0_clk,                 --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,      -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,    --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,     --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,    --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,   --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,    --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,   --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,    --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,   --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,   --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,       --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,     --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,     --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,     --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,    --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,    --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,       --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,     --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,    --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,    --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,      --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,    --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,     --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,    --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,   --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,    --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,   --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,    --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,   --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,   --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,       --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,     --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,     --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,     --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,    --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready     --                  .rready
		);

	jtag_uart_0 : component soc_system_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver1_irq                                     --               irq.irq
		);

	matches_mutex : component soc_system_finished_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,      -- reset.reset_n
			clk           => pll_0_outclk0_clk,                             --   clk.clk
			chipselect    => mm_interconnect_0_matches_mutex_s1_chipselect, --    s1.chipselect
			data_from_cpu => mm_interconnect_0_matches_mutex_s1_writedata,  --      .writedata
			read          => mm_interconnect_0_matches_mutex_s1_read,       --      .read
			write         => mm_interconnect_0_matches_mutex_s1_write,      --      .write
			data_to_cpu   => mm_interconnect_0_matches_mutex_s1_readdata,   --      .readdata
			address       => mm_interconnect_0_matches_mutex_s1_address(0)  --      .address
		);

	paper_mutex : component soc_system_finished_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,    -- reset.reset_n
			clk           => pll_0_outclk0_clk,                           --   clk.clk
			chipselect    => mm_interconnect_0_paper_mutex_s1_chipselect, --    s1.chipselect
			data_from_cpu => mm_interconnect_0_paper_mutex_s1_writedata,  --      .writedata
			read          => mm_interconnect_0_paper_mutex_s1_read,       --      .read
			write         => mm_interconnect_0_paper_mutex_s1_write,      --      .write
			data_to_cpu   => mm_interconnect_0_paper_mutex_s1_readdata,   --      .readdata
			address       => mm_interconnect_0_paper_mutex_s1_address(0)  --      .address
		);

	pll_0 : component soc_system_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			outclk_1 => pll_0_outclk1_clk,       -- outclk1.clk
			outclk_2 => pll_0_sdram_clk,         -- outclk2.clk
			locked   => open                     -- (terminated)
		);

	sdram_controller_0 : component soc_system_sdram_controller_0
		port map (
			clk            => pll_0_outclk1_clk,                                            --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,                 -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_0_wire_we_n                                  --      .export
		);

	smoker_with_matches : component soc_system_smoker_with_matches
		port map (
			clk                                 => clk_clk,                                                           --                       clk.clk
			reset_n                             => rst_controller_003_reset_out_reset_ports_inv,                      --                     reset.reset_n
			reset_req                           => rst_controller_003_reset_out_reset_req,                            --                          .reset_req
			d_address                           => smoker_with_matches_data_master_address,                           --               data_master.address
			d_byteenable                        => smoker_with_matches_data_master_byteenable,                        --                          .byteenable
			d_read                              => smoker_with_matches_data_master_read,                              --                          .read
			d_readdata                          => smoker_with_matches_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => smoker_with_matches_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => smoker_with_matches_data_master_write,                             --                          .write
			d_writedata                         => smoker_with_matches_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => smoker_with_matches_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => smoker_with_matches_instruction_master_address,                    --        instruction_master.address
			i_read                              => smoker_with_matches_instruction_master_read,                       --                          .read
			i_readdata                          => smoker_with_matches_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => smoker_with_matches_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => smoker_with_matches_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => smoker_with_matches_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_smoker_with_matches_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_smoker_with_matches_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_smoker_with_matches_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_smoker_with_matches_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_smoker_with_matches_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_smoker_with_matches_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_smoker_with_matches_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_smoker_with_matches_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                               -- custom_instruction_master.readra
		);

	smoker_with_paper : component soc_system_smoker_with_paper
		port map (
			clk                                 => pll_0_outclk0_clk,                                               --                       clk.clk
			reset_n                             => rst_controller_004_reset_out_reset_ports_inv,                    --                     reset.reset_n
			reset_req                           => rst_controller_004_reset_out_reset_req,                          --                          .reset_req
			d_address                           => smoker_with_paper_data_master_address,                           --               data_master.address
			d_byteenable                        => smoker_with_paper_data_master_byteenable,                        --                          .byteenable
			d_read                              => smoker_with_paper_data_master_read,                              --                          .read
			d_readdata                          => smoker_with_paper_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => smoker_with_paper_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => smoker_with_paper_data_master_write,                             --                          .write
			d_writedata                         => smoker_with_paper_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => smoker_with_paper_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => smoker_with_paper_instruction_master_address,                    --        instruction_master.address
			i_read                              => smoker_with_paper_instruction_master_read,                       --                          .read
			i_readdata                          => smoker_with_paper_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => smoker_with_paper_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => smoker_with_paper_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => smoker_with_paper_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_smoker_with_paper_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_smoker_with_paper_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_smoker_with_paper_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_smoker_with_paper_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_smoker_with_paper_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_smoker_with_paper_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_smoker_with_paper_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_smoker_with_paper_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                             -- custom_instruction_master.readra
		);

	smoker_with_tobacco : component soc_system_smoker_with_tobacco
		port map (
			clk                                 => pll_0_outclk0_clk,                                                 --                       clk.clk
			reset_n                             => rst_controller_005_reset_out_reset_ports_inv,                      --                     reset.reset_n
			reset_req                           => rst_controller_005_reset_out_reset_req,                            --                          .reset_req
			d_address                           => smoker_with_tobacco_data_master_address,                           --               data_master.address
			d_byteenable                        => smoker_with_tobacco_data_master_byteenable,                        --                          .byteenable
			d_read                              => smoker_with_tobacco_data_master_read,                              --                          .read
			d_readdata                          => smoker_with_tobacco_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => smoker_with_tobacco_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => smoker_with_tobacco_data_master_write,                             --                          .write
			d_writedata                         => smoker_with_tobacco_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => smoker_with_tobacco_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => smoker_with_tobacco_instruction_master_address,                    --        instruction_master.address
			i_read                              => smoker_with_tobacco_instruction_master_read,                       --                          .read
			i_readdata                          => smoker_with_tobacco_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => smoker_with_tobacco_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => smoker_with_tobacco_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => smoker_with_tobacco_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                               -- custom_instruction_master.readra
		);

	sysid : component soc_system_sysid
		port map (
			clock    => pll_0_outclk0_clk,                                --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_0 : component soc_system_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_005_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_002_receiver1_irq                  --   irq.irq
		);

	timer_1 : component soc_system_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_006_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_001_receiver0_irq                  --   irq.irq
		);

	timer_2 : component soc_system_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_007_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_2_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_2_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_2_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_2_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_2_s1_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_receiver_irq(0)              --   irq.irq
		);

	tobacco_mutex : component soc_system_finished_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,      -- reset.reset_n
			clk           => pll_0_outclk0_clk,                             --   clk.clk
			chipselect    => mm_interconnect_0_tobacco_mutex_s1_chipselect, --    s1.chipselect
			data_from_cpu => mm_interconnect_0_tobacco_mutex_s1_writedata,  --      .writedata
			read          => mm_interconnect_0_tobacco_mutex_s1_read,       --      .read
			write         => mm_interconnect_0_tobacco_mutex_s1_write,      --      .write
			data_to_cpu   => mm_interconnect_0_tobacco_mutex_s1_readdata,   --      .readdata
			address       => mm_interconnect_0_tobacco_mutex_s1_address(0)  --      .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                      --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                                    --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                     --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                                    --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                                   --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                                    --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                                   --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                                    --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                                   --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                                   --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                       --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                     --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                     --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                     --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                                    --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                                    --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                       --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                     --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                                    --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                                    --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                      --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                                    --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                     --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                                    --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                                   --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                                    --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                                   --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                                    --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                                   --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                                   --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                       --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                     --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                     --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                     --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                                    --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                                    --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                           --                                                     clk_0_clk.clk
			pll_0_outclk0_clk                                                   => pll_0_outclk0_clk,                                                 --                                                 pll_0_outclk0.clk
			pll_0_outclk1_clk                                                   => pll_0_outclk1_clk,                                                 --                                                 pll_0_outclk1.clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_008_reset_out_reset,                                -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset                       => rst_controller_001_reset_out_reset,                                --                       jtag_uart_0_reset_reset_bridge_in_reset.reset
			sdram_controller_0_reset_reset_bridge_in_reset_reset                => rst_controller_002_reset_out_reset,                                --                sdram_controller_0_reset_reset_bridge_in_reset.reset
			smoker_with_matches_reset_reset_bridge_in_reset_reset               => rst_controller_003_reset_out_reset,                                --               smoker_with_matches_reset_reset_bridge_in_reset.reset
			smoker_with_paper_reset_reset_bridge_in_reset_reset                 => rst_controller_004_reset_out_reset,                                --                 smoker_with_paper_reset_reset_bridge_in_reset.reset
			smoker_with_tobacco_reset_reset_bridge_in_reset_reset               => rst_controller_005_reset_out_reset,                                --               smoker_with_tobacco_reset_reset_bridge_in_reset.reset
			timer_1_reset_reset_bridge_in_reset_reset                           => rst_controller_006_reset_out_reset,                                --                           timer_1_reset_reset_bridge_in_reset.reset
			timer_2_reset_reset_bridge_in_reset_reset                           => rst_controller_007_reset_out_reset,                                --                           timer_2_reset_reset_bridge_in_reset.reset
			tobacco_mutex_reset_reset_bridge_in_reset_reset                     => rst_controller_reset_out_reset,                                    --                     tobacco_mutex_reset_reset_bridge_in_reset.reset
			smoker_with_matches_data_master_address                             => smoker_with_matches_data_master_address,                           --                               smoker_with_matches_data_master.address
			smoker_with_matches_data_master_waitrequest                         => smoker_with_matches_data_master_waitrequest,                       --                                                              .waitrequest
			smoker_with_matches_data_master_byteenable                          => smoker_with_matches_data_master_byteenable,                        --                                                              .byteenable
			smoker_with_matches_data_master_read                                => smoker_with_matches_data_master_read,                              --                                                              .read
			smoker_with_matches_data_master_readdata                            => smoker_with_matches_data_master_readdata,                          --                                                              .readdata
			smoker_with_matches_data_master_write                               => smoker_with_matches_data_master_write,                             --                                                              .write
			smoker_with_matches_data_master_writedata                           => smoker_with_matches_data_master_writedata,                         --                                                              .writedata
			smoker_with_matches_data_master_debugaccess                         => smoker_with_matches_data_master_debugaccess,                       --                                                              .debugaccess
			smoker_with_matches_instruction_master_address                      => smoker_with_matches_instruction_master_address,                    --                        smoker_with_matches_instruction_master.address
			smoker_with_matches_instruction_master_waitrequest                  => smoker_with_matches_instruction_master_waitrequest,                --                                                              .waitrequest
			smoker_with_matches_instruction_master_read                         => smoker_with_matches_instruction_master_read,                       --                                                              .read
			smoker_with_matches_instruction_master_readdata                     => smoker_with_matches_instruction_master_readdata,                   --                                                              .readdata
			smoker_with_paper_data_master_address                               => smoker_with_paper_data_master_address,                             --                                 smoker_with_paper_data_master.address
			smoker_with_paper_data_master_waitrequest                           => smoker_with_paper_data_master_waitrequest,                         --                                                              .waitrequest
			smoker_with_paper_data_master_byteenable                            => smoker_with_paper_data_master_byteenable,                          --                                                              .byteenable
			smoker_with_paper_data_master_read                                  => smoker_with_paper_data_master_read,                                --                                                              .read
			smoker_with_paper_data_master_readdata                              => smoker_with_paper_data_master_readdata,                            --                                                              .readdata
			smoker_with_paper_data_master_write                                 => smoker_with_paper_data_master_write,                               --                                                              .write
			smoker_with_paper_data_master_writedata                             => smoker_with_paper_data_master_writedata,                           --                                                              .writedata
			smoker_with_paper_data_master_debugaccess                           => smoker_with_paper_data_master_debugaccess,                         --                                                              .debugaccess
			smoker_with_paper_instruction_master_address                        => smoker_with_paper_instruction_master_address,                      --                          smoker_with_paper_instruction_master.address
			smoker_with_paper_instruction_master_waitrequest                    => smoker_with_paper_instruction_master_waitrequest,                  --                                                              .waitrequest
			smoker_with_paper_instruction_master_read                           => smoker_with_paper_instruction_master_read,                         --                                                              .read
			smoker_with_paper_instruction_master_readdata                       => smoker_with_paper_instruction_master_readdata,                     --                                                              .readdata
			smoker_with_tobacco_data_master_address                             => smoker_with_tobacco_data_master_address,                           --                               smoker_with_tobacco_data_master.address
			smoker_with_tobacco_data_master_waitrequest                         => smoker_with_tobacco_data_master_waitrequest,                       --                                                              .waitrequest
			smoker_with_tobacco_data_master_byteenable                          => smoker_with_tobacco_data_master_byteenable,                        --                                                              .byteenable
			smoker_with_tobacco_data_master_read                                => smoker_with_tobacco_data_master_read,                              --                                                              .read
			smoker_with_tobacco_data_master_readdata                            => smoker_with_tobacco_data_master_readdata,                          --                                                              .readdata
			smoker_with_tobacco_data_master_write                               => smoker_with_tobacco_data_master_write,                             --                                                              .write
			smoker_with_tobacco_data_master_writedata                           => smoker_with_tobacco_data_master_writedata,                         --                                                              .writedata
			smoker_with_tobacco_data_master_debugaccess                         => smoker_with_tobacco_data_master_debugaccess,                       --                                                              .debugaccess
			smoker_with_tobacco_instruction_master_address                      => smoker_with_tobacco_instruction_master_address,                    --                        smoker_with_tobacco_instruction_master.address
			smoker_with_tobacco_instruction_master_waitrequest                  => smoker_with_tobacco_instruction_master_waitrequest,                --                                                              .waitrequest
			smoker_with_tobacco_instruction_master_read                         => smoker_with_tobacco_instruction_master_read,                       --                                                              .read
			smoker_with_tobacco_instruction_master_readdata                     => smoker_with_tobacco_instruction_master_readdata,                   --                                                              .readdata
			finished_mutex_s1_address                                           => mm_interconnect_0_finished_mutex_s1_address,                       --                                             finished_mutex_s1.address
			finished_mutex_s1_write                                             => mm_interconnect_0_finished_mutex_s1_write,                         --                                                              .write
			finished_mutex_s1_read                                              => mm_interconnect_0_finished_mutex_s1_read,                          --                                                              .read
			finished_mutex_s1_readdata                                          => mm_interconnect_0_finished_mutex_s1_readdata,                      --                                                              .readdata
			finished_mutex_s1_writedata                                         => mm_interconnect_0_finished_mutex_s1_writedata,                     --                                                              .writedata
			finished_mutex_s1_chipselect                                        => mm_interconnect_0_finished_mutex_s1_chipselect,                    --                                                              .chipselect
			jtag_uart_0_avalon_jtag_slave_address                               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,           --                                 jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,             --                                                              .write
			jtag_uart_0_avalon_jtag_slave_read                                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,              --                                                              .read
			jtag_uart_0_avalon_jtag_slave_readdata                              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,          --                                                              .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,         --                                                              .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,       --                                                              .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,        --                                                              .chipselect
			matches_mutex_s1_address                                            => mm_interconnect_0_matches_mutex_s1_address,                        --                                              matches_mutex_s1.address
			matches_mutex_s1_write                                              => mm_interconnect_0_matches_mutex_s1_write,                          --                                                              .write
			matches_mutex_s1_read                                               => mm_interconnect_0_matches_mutex_s1_read,                           --                                                              .read
			matches_mutex_s1_readdata                                           => mm_interconnect_0_matches_mutex_s1_readdata,                       --                                                              .readdata
			matches_mutex_s1_writedata                                          => mm_interconnect_0_matches_mutex_s1_writedata,                      --                                                              .writedata
			matches_mutex_s1_chipselect                                         => mm_interconnect_0_matches_mutex_s1_chipselect,                     --                                                              .chipselect
			paper_mutex_s1_address                                              => mm_interconnect_0_paper_mutex_s1_address,                          --                                                paper_mutex_s1.address
			paper_mutex_s1_write                                                => mm_interconnect_0_paper_mutex_s1_write,                            --                                                              .write
			paper_mutex_s1_read                                                 => mm_interconnect_0_paper_mutex_s1_read,                             --                                                              .read
			paper_mutex_s1_readdata                                             => mm_interconnect_0_paper_mutex_s1_readdata,                         --                                                              .readdata
			paper_mutex_s1_writedata                                            => mm_interconnect_0_paper_mutex_s1_writedata,                        --                                                              .writedata
			paper_mutex_s1_chipselect                                           => mm_interconnect_0_paper_mutex_s1_chipselect,                       --                                                              .chipselect
			sdram_controller_0_s1_address                                       => mm_interconnect_0_sdram_controller_0_s1_address,                   --                                         sdram_controller_0_s1.address
			sdram_controller_0_s1_write                                         => mm_interconnect_0_sdram_controller_0_s1_write,                     --                                                              .write
			sdram_controller_0_s1_read                                          => mm_interconnect_0_sdram_controller_0_s1_read,                      --                                                              .read
			sdram_controller_0_s1_readdata                                      => mm_interconnect_0_sdram_controller_0_s1_readdata,                  --                                                              .readdata
			sdram_controller_0_s1_writedata                                     => mm_interconnect_0_sdram_controller_0_s1_writedata,                 --                                                              .writedata
			sdram_controller_0_s1_byteenable                                    => mm_interconnect_0_sdram_controller_0_s1_byteenable,                --                                                              .byteenable
			sdram_controller_0_s1_readdatavalid                                 => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,             --                                                              .readdatavalid
			sdram_controller_0_s1_waitrequest                                   => mm_interconnect_0_sdram_controller_0_s1_waitrequest,               --                                                              .waitrequest
			sdram_controller_0_s1_chipselect                                    => mm_interconnect_0_sdram_controller_0_s1_chipselect,                --                                                              .chipselect
			smoker_with_matches_debug_mem_slave_address                         => mm_interconnect_0_smoker_with_matches_debug_mem_slave_address,     --                           smoker_with_matches_debug_mem_slave.address
			smoker_with_matches_debug_mem_slave_write                           => mm_interconnect_0_smoker_with_matches_debug_mem_slave_write,       --                                                              .write
			smoker_with_matches_debug_mem_slave_read                            => mm_interconnect_0_smoker_with_matches_debug_mem_slave_read,        --                                                              .read
			smoker_with_matches_debug_mem_slave_readdata                        => mm_interconnect_0_smoker_with_matches_debug_mem_slave_readdata,    --                                                              .readdata
			smoker_with_matches_debug_mem_slave_writedata                       => mm_interconnect_0_smoker_with_matches_debug_mem_slave_writedata,   --                                                              .writedata
			smoker_with_matches_debug_mem_slave_byteenable                      => mm_interconnect_0_smoker_with_matches_debug_mem_slave_byteenable,  --                                                              .byteenable
			smoker_with_matches_debug_mem_slave_waitrequest                     => mm_interconnect_0_smoker_with_matches_debug_mem_slave_waitrequest, --                                                              .waitrequest
			smoker_with_matches_debug_mem_slave_debugaccess                     => mm_interconnect_0_smoker_with_matches_debug_mem_slave_debugaccess, --                                                              .debugaccess
			smoker_with_paper_debug_mem_slave_address                           => mm_interconnect_0_smoker_with_paper_debug_mem_slave_address,       --                             smoker_with_paper_debug_mem_slave.address
			smoker_with_paper_debug_mem_slave_write                             => mm_interconnect_0_smoker_with_paper_debug_mem_slave_write,         --                                                              .write
			smoker_with_paper_debug_mem_slave_read                              => mm_interconnect_0_smoker_with_paper_debug_mem_slave_read,          --                                                              .read
			smoker_with_paper_debug_mem_slave_readdata                          => mm_interconnect_0_smoker_with_paper_debug_mem_slave_readdata,      --                                                              .readdata
			smoker_with_paper_debug_mem_slave_writedata                         => mm_interconnect_0_smoker_with_paper_debug_mem_slave_writedata,     --                                                              .writedata
			smoker_with_paper_debug_mem_slave_byteenable                        => mm_interconnect_0_smoker_with_paper_debug_mem_slave_byteenable,    --                                                              .byteenable
			smoker_with_paper_debug_mem_slave_waitrequest                       => mm_interconnect_0_smoker_with_paper_debug_mem_slave_waitrequest,   --                                                              .waitrequest
			smoker_with_paper_debug_mem_slave_debugaccess                       => mm_interconnect_0_smoker_with_paper_debug_mem_slave_debugaccess,   --                                                              .debugaccess
			smoker_with_tobacco_debug_mem_slave_address                         => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_address,     --                           smoker_with_tobacco_debug_mem_slave.address
			smoker_with_tobacco_debug_mem_slave_write                           => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_write,       --                                                              .write
			smoker_with_tobacco_debug_mem_slave_read                            => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_read,        --                                                              .read
			smoker_with_tobacco_debug_mem_slave_readdata                        => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_readdata,    --                                                              .readdata
			smoker_with_tobacco_debug_mem_slave_writedata                       => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_writedata,   --                                                              .writedata
			smoker_with_tobacco_debug_mem_slave_byteenable                      => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_byteenable,  --                                                              .byteenable
			smoker_with_tobacco_debug_mem_slave_waitrequest                     => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_waitrequest, --                                                              .waitrequest
			smoker_with_tobacco_debug_mem_slave_debugaccess                     => mm_interconnect_0_smoker_with_tobacco_debug_mem_slave_debugaccess, --                                                              .debugaccess
			sysid_control_slave_address                                         => mm_interconnect_0_sysid_control_slave_address,                     --                                           sysid_control_slave.address
			sysid_control_slave_readdata                                        => mm_interconnect_0_sysid_control_slave_readdata,                    --                                                              .readdata
			timer_0_s1_address                                                  => mm_interconnect_0_timer_0_s1_address,                              --                                                    timer_0_s1.address
			timer_0_s1_write                                                    => mm_interconnect_0_timer_0_s1_write,                                --                                                              .write
			timer_0_s1_readdata                                                 => mm_interconnect_0_timer_0_s1_readdata,                             --                                                              .readdata
			timer_0_s1_writedata                                                => mm_interconnect_0_timer_0_s1_writedata,                            --                                                              .writedata
			timer_0_s1_chipselect                                               => mm_interconnect_0_timer_0_s1_chipselect,                           --                                                              .chipselect
			timer_1_s1_address                                                  => mm_interconnect_0_timer_1_s1_address,                              --                                                    timer_1_s1.address
			timer_1_s1_write                                                    => mm_interconnect_0_timer_1_s1_write,                                --                                                              .write
			timer_1_s1_readdata                                                 => mm_interconnect_0_timer_1_s1_readdata,                             --                                                              .readdata
			timer_1_s1_writedata                                                => mm_interconnect_0_timer_1_s1_writedata,                            --                                                              .writedata
			timer_1_s1_chipselect                                               => mm_interconnect_0_timer_1_s1_chipselect,                           --                                                              .chipselect
			timer_2_s1_address                                                  => mm_interconnect_0_timer_2_s1_address,                              --                                                    timer_2_s1.address
			timer_2_s1_write                                                    => mm_interconnect_0_timer_2_s1_write,                                --                                                              .write
			timer_2_s1_readdata                                                 => mm_interconnect_0_timer_2_s1_readdata,                             --                                                              .readdata
			timer_2_s1_writedata                                                => mm_interconnect_0_timer_2_s1_writedata,                            --                                                              .writedata
			timer_2_s1_chipselect                                               => mm_interconnect_0_timer_2_s1_chipselect,                           --                                                              .chipselect
			tobacco_mutex_s1_address                                            => mm_interconnect_0_tobacco_mutex_s1_address,                        --                                              tobacco_mutex_s1.address
			tobacco_mutex_s1_write                                              => mm_interconnect_0_tobacco_mutex_s1_write,                          --                                                              .write
			tobacco_mutex_s1_read                                               => mm_interconnect_0_tobacco_mutex_s1_read,                           --                                                              .read
			tobacco_mutex_s1_readdata                                           => mm_interconnect_0_tobacco_mutex_s1_readdata,                       --                                                              .readdata
			tobacco_mutex_s1_writedata                                          => mm_interconnect_0_tobacco_mutex_s1_writedata,                      --                                                              .writedata
			tobacco_mutex_s1_chipselect                                         => mm_interconnect_0_tobacco_mutex_s1_chipselect                      --                                                              .chipselect
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_003_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => smoker_with_matches_irq_irq         --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,                  --       clk.clk
			reset         => rst_controller_004_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_001_receiver1_irq,       -- receiver1.irq
			sender_irq    => smoker_with_paper_irq_irq           --    sender.irq
		);

	irq_mapper_002 : component soc_system_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,                  --       clk.clk
			reset         => rst_controller_005_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver1_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_002_receiver1_irq,       -- receiver1.irq
			sender_irq    => smoker_with_tobacco_irq_irq         --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => clk_clk,                            --         sender_clk.clk
			receiver_reset => rst_controller_007_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_003_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk    => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk      => clk_clk,                            --         sender_clk.clk
			receiver_reset  => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset    => rst_controller_003_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq(0) => irq_mapper_001_receiver1_irq,       --           receiver.irq
			sender_irq(0)   => irq_mapper_receiver1_irq            --             sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                       -- reset_in0.reset
			reset_in1      => smoker_with_tobacco_debug_reset_request_reset, -- reset_in1.reset
			reset_in2      => smoker_with_paper_debug_reset_request_reset,   -- reset_in2.reset
			clk            => pll_0_outclk0_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,                -- reset_out.reset
			reset_req      => open,                                          -- (terminated)
			reset_req_in0  => '0',                                           -- (terminated)
			reset_req_in1  => '0',                                           -- (terminated)
			reset_req_in2  => '0',                                           -- (terminated)
			reset_in3      => '0',                                           -- (terminated)
			reset_req_in3  => '0',                                           -- (terminated)
			reset_in4      => '0',                                           -- (terminated)
			reset_req_in4  => '0',                                           -- (terminated)
			reset_in5      => '0',                                           -- (terminated)
			reset_req_in5  => '0',                                           -- (terminated)
			reset_in6      => '0',                                           -- (terminated)
			reset_req_in6  => '0',                                           -- (terminated)
			reset_in7      => '0',                                           -- (terminated)
			reset_req_in7  => '0',                                           -- (terminated)
			reset_in8      => '0',                                           -- (terminated)
			reset_req_in8  => '0',                                           -- (terminated)
			reset_in9      => '0',                                           -- (terminated)
			reset_req_in9  => '0',                                           -- (terminated)
			reset_in10     => '0',                                           -- (terminated)
			reset_req_in10 => '0',                                           -- (terminated)
			reset_in11     => '0',                                           -- (terminated)
			reset_req_in11 => '0',                                           -- (terminated)
			reset_in12     => '0',                                           -- (terminated)
			reset_req_in12 => '0',                                           -- (terminated)
			reset_in13     => '0',                                           -- (terminated)
			reset_req_in13 => '0',                                           -- (terminated)
			reset_in14     => '0',                                           -- (terminated)
			reset_req_in14 => '0',                                           -- (terminated)
			reset_in15     => '0',                                           -- (terminated)
			reset_req_in15 => '0'                                            -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 4,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                       -- reset_in0.reset
			reset_in1      => smoker_with_tobacco_debug_reset_request_reset, -- reset_in1.reset
			reset_in2      => smoker_with_paper_debug_reset_request_reset,   -- reset_in2.reset
			reset_in3      => smoker_with_matches_debug_reset_request_reset, -- reset_in3.reset
			clk            => pll_0_outclk0_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,            -- reset_out.reset
			reset_req      => open,                                          -- (terminated)
			reset_req_in0  => '0',                                           -- (terminated)
			reset_req_in1  => '0',                                           -- (terminated)
			reset_req_in2  => '0',                                           -- (terminated)
			reset_req_in3  => '0',                                           -- (terminated)
			reset_in4      => '0',                                           -- (terminated)
			reset_req_in4  => '0',                                           -- (terminated)
			reset_in5      => '0',                                           -- (terminated)
			reset_req_in5  => '0',                                           -- (terminated)
			reset_in6      => '0',                                           -- (terminated)
			reset_req_in6  => '0',                                           -- (terminated)
			reset_in7      => '0',                                           -- (terminated)
			reset_req_in7  => '0',                                           -- (terminated)
			reset_in8      => '0',                                           -- (terminated)
			reset_req_in8  => '0',                                           -- (terminated)
			reset_in9      => '0',                                           -- (terminated)
			reset_req_in9  => '0',                                           -- (terminated)
			reset_in10     => '0',                                           -- (terminated)
			reset_req_in10 => '0',                                           -- (terminated)
			reset_in11     => '0',                                           -- (terminated)
			reset_req_in11 => '0',                                           -- (terminated)
			reset_in12     => '0',                                           -- (terminated)
			reset_req_in12 => '0',                                           -- (terminated)
			reset_in13     => '0',                                           -- (terminated)
			reset_req_in13 => '0',                                           -- (terminated)
			reset_in14     => '0',                                           -- (terminated)
			reset_req_in14 => '0',                                           -- (terminated)
			reset_in15     => '0',                                           -- (terminated)
			reset_req_in15 => '0'                                            -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_0_outclk1_clk,                  --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component soc_system_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_003_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_004 : component soc_system_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_004_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_005 : component soc_system_rst_controller_005
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                       -- reset_in0.reset
			reset_in1      => smoker_with_tobacco_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                             --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset,            -- reset_out.reset
			reset_req      => rst_controller_005_reset_out_reset_req,        --          .reset_req
			reset_req_in0  => '0',                                           -- (terminated)
			reset_req_in1  => '0',                                           -- (terminated)
			reset_in2      => '0',                                           -- (terminated)
			reset_req_in2  => '0',                                           -- (terminated)
			reset_in3      => '0',                                           -- (terminated)
			reset_req_in3  => '0',                                           -- (terminated)
			reset_in4      => '0',                                           -- (terminated)
			reset_req_in4  => '0',                                           -- (terminated)
			reset_in5      => '0',                                           -- (terminated)
			reset_req_in5  => '0',                                           -- (terminated)
			reset_in6      => '0',                                           -- (terminated)
			reset_req_in6  => '0',                                           -- (terminated)
			reset_in7      => '0',                                           -- (terminated)
			reset_req_in7  => '0',                                           -- (terminated)
			reset_in8      => '0',                                           -- (terminated)
			reset_req_in8  => '0',                                           -- (terminated)
			reset_in9      => '0',                                           -- (terminated)
			reset_req_in9  => '0',                                           -- (terminated)
			reset_in10     => '0',                                           -- (terminated)
			reset_req_in10 => '0',                                           -- (terminated)
			reset_in11     => '0',                                           -- (terminated)
			reset_req_in11 => '0',                                           -- (terminated)
			reset_in12     => '0',                                           -- (terminated)
			reset_req_in12 => '0',                                           -- (terminated)
			reset_in13     => '0',                                           -- (terminated)
			reset_req_in13 => '0',                                           -- (terminated)
			reset_in14     => '0',                                           -- (terminated)
			reset_req_in14 => '0',                                           -- (terminated)
			reset_in15     => '0',                                           -- (terminated)
			reset_req_in15 => '0'                                            -- (terminated)
		);

	rst_controller_006 : component soc_system_rst_controller_006
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                     -- reset_in0.reset
			reset_in1      => smoker_with_paper_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                           --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset,          -- reset_out.reset
			reset_req      => open,                                        -- (terminated)
			reset_req_in0  => '0',                                         -- (terminated)
			reset_req_in1  => '0',                                         -- (terminated)
			reset_in2      => '0',                                         -- (terminated)
			reset_req_in2  => '0',                                         -- (terminated)
			reset_in3      => '0',                                         -- (terminated)
			reset_req_in3  => '0',                                         -- (terminated)
			reset_in4      => '0',                                         -- (terminated)
			reset_req_in4  => '0',                                         -- (terminated)
			reset_in5      => '0',                                         -- (terminated)
			reset_req_in5  => '0',                                         -- (terminated)
			reset_in6      => '0',                                         -- (terminated)
			reset_req_in6  => '0',                                         -- (terminated)
			reset_in7      => '0',                                         -- (terminated)
			reset_req_in7  => '0',                                         -- (terminated)
			reset_in8      => '0',                                         -- (terminated)
			reset_req_in8  => '0',                                         -- (terminated)
			reset_in9      => '0',                                         -- (terminated)
			reset_req_in9  => '0',                                         -- (terminated)
			reset_in10     => '0',                                         -- (terminated)
			reset_req_in10 => '0',                                         -- (terminated)
			reset_in11     => '0',                                         -- (terminated)
			reset_req_in11 => '0',                                         -- (terminated)
			reset_in12     => '0',                                         -- (terminated)
			reset_req_in12 => '0',                                         -- (terminated)
			reset_in13     => '0',                                         -- (terminated)
			reset_req_in13 => '0',                                         -- (terminated)
			reset_in14     => '0',                                         -- (terminated)
			reset_req_in14 => '0',                                         -- (terminated)
			reset_in15     => '0',                                         -- (terminated)
			reset_req_in15 => '0'                                          -- (terminated)
		);

	rst_controller_007 : component soc_system_rst_controller_006
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                       -- reset_in0.reset
			reset_in1      => smoker_with_matches_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                             --       clk.clk
			reset_out      => rst_controller_007_reset_out_reset,            -- reset_out.reset
			reset_req      => open,                                          -- (terminated)
			reset_req_in0  => '0',                                           -- (terminated)
			reset_req_in1  => '0',                                           -- (terminated)
			reset_in2      => '0',                                           -- (terminated)
			reset_req_in2  => '0',                                           -- (terminated)
			reset_in3      => '0',                                           -- (terminated)
			reset_req_in3  => '0',                                           -- (terminated)
			reset_in4      => '0',                                           -- (terminated)
			reset_req_in4  => '0',                                           -- (terminated)
			reset_in5      => '0',                                           -- (terminated)
			reset_req_in5  => '0',                                           -- (terminated)
			reset_in6      => '0',                                           -- (terminated)
			reset_req_in6  => '0',                                           -- (terminated)
			reset_in7      => '0',                                           -- (terminated)
			reset_req_in7  => '0',                                           -- (terminated)
			reset_in8      => '0',                                           -- (terminated)
			reset_req_in8  => '0',                                           -- (terminated)
			reset_in9      => '0',                                           -- (terminated)
			reset_req_in9  => '0',                                           -- (terminated)
			reset_in10     => '0',                                           -- (terminated)
			reset_req_in10 => '0',                                           -- (terminated)
			reset_in11     => '0',                                           -- (terminated)
			reset_req_in11 => '0',                                           -- (terminated)
			reset_in12     => '0',                                           -- (terminated)
			reset_req_in12 => '0',                                           -- (terminated)
			reset_in13     => '0',                                           -- (terminated)
			reset_req_in13 => '0',                                           -- (terminated)
			reset_in14     => '0',                                           -- (terminated)
			reset_req_in14 => '0',                                           -- (terminated)
			reset_in15     => '0',                                           -- (terminated)
			reset_req_in15 => '0'                                            -- (terminated)
		);

	rst_controller_008 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_008_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	mm_interconnect_0_timer_2_s1_write_ports_inv <= not mm_interconnect_0_timer_2_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	rst_controller_005_reset_out_reset_ports_inv <= not rst_controller_005_reset_out_reset;

	rst_controller_006_reset_out_reset_ports_inv <= not rst_controller_006_reset_out_reset;

	rst_controller_007_reset_out_reset_ports_inv <= not rst_controller_007_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system
