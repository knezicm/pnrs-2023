
module soc_system (
	clk_clk,
	leds_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output	[9:0]	leds_0_external_connection_export;
	input		reset_reset_n;
endmodule
